module q4(m,p,q);
input [2:0]m,q;
output [3:0]p;
wire [3:1]c1,c2;
assign p[0]=m[0] & q[0];
assign p[1]=fa ;

