`timescale 1ns/1ns
`include "mux16.v"

module mux16_tb;
reg [3:0]s;
reg[15:0]w;
wire f;
mux16 vvt(s,w,f);
initial begin
 
 $dumpfile("mux16_tb.vcd");
 $dumpvars(0,mux16_tb);

s=0; 
w=16'b1110000111000001;
#20
 
 s=1; 
w=16'b1110000111000001;
#20
 
 s=2; 
w=16'b1110000111000001;
#20
 
 s=3; 
w=16'b1110000111000001;
#20
 
 s=4; 
w=16'b1110000111000001;
#20
 
 s=5; 
w=16'b1110000111000001;
#20
 
 s=6; 
w=16'b1110000111000001;
#20
 
 s=7; 
w=16'b1110000111000001;
#20
 
 s=8; 
w=16'b1110000111000001;
#20
 
 s=9; 
w=16'b1110000111000001;
#20
 
 s=10; 
w=16'b1110000111000001;
#20
 
 s=11; 
w=16'b1110000111000001;
#20
 
 s=12; 
w=16'b1110000111000001;
#20
 
 s=13; 
w=16'b1110000111000001;
#20
 
 s=14; 
w=16'b1110000111000001;
#20
 
 s=15; 
w=16'b1110000111000001;
#20
 
$display("Test complete");
 end
 endmodule
